///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
///////////////////////////////////////////

    Zihpm_cg = new();    Zihpm_cg.set_inst_name("obj_Zihpm");