///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
///////////////////////////////////////////

`define COVER_ZIHPM
covergroup Zihpm_cg with function sample (ins_t, ins);
    option.per_instance = 0;
    `include "coverage/RISCV_coverage_standard_coverpoints.svh"

cp_hpm_count: coverpoint {ins.current.insn[31:20], ins.current.csr[12'hB03][31:0] } {
        bins cycle_enabled         = {44'b110000000000_00000000000000000000000000000001};
        bins time_enabled          = {44'b110000000001_00000000000000000000000000000010};
        bins instret_enabled       = {44'b110000000010_00000000000000000000000000000100};
        bins mhpmcounter3_enabled   = {44'b110000000011_00000000000000000000000000001000};
        bins mhpmcounter4_enabled   = {44'b110000000100_00000000000000000000000000010000};
        bins mhpmcounter5_enabled   = {44'b110000000101_00000000000000000000000000100000};
        bins mhpmcounter6_enabled   = {44'b110000000110_00000000000000000000000001000000};
        bins mhpmcounter7_enabled   = {44'b110000000111_00000000000000000000000010000000};
        bins mhpmcounter8_enabled   = {44'b110000001000_00000000000000000000000100000000};
        bins mhpmcounter9_enabled   = {44'b110000001001_00000000000000000000001000000000};
        bins mhpmcounter10_enabled  = {44'b110000001010_00000000000000000000010000000000};
        bins mhpmcounter11_enabled  = {44'b110000001011_00000000000000000000100000000000};
        bins mhpmcounter12_enabled  = {44'b110000001100_00000000000000000001000000000000};
        bins mhpmcounter13_enabled  = {44'b110000001101_00000000000000000010000000000000};
        bins mhpmcounter14_enabled  = {44'b110000001110_00000000000000000100000000000000};
        bins mhpmcounter15_enabled  = {44'b110000001111_00000000000000001000000000000000};
        bins mhpmcounter16_enabled  = {44'b110000010000_00000000000000010000000000000000};
        bins mhpmcounter17_enabled  = {44'b110000010001_00000000000000100000000000000000};
        bins mhpmcounter18_enabled  = {44'b110000010010_00000000000001000000000000000000};
        bins mhpmcounter19_enabled  = {44'b110000010011_00000000000010000000000000000000};
        bins mhpmcounter20_enabled  = {44'b110000010100_00000000000100000000000000000000};
        bins mhpmcounter21_enabled  = {44'b110000010101_00000000001000000000000000000000};
        bins mhpmcounter22_enabled  = {44'b110000010110_00000000010000000000000000000000};
        bins mhpmcounter23_enabled  = {44'b110000010111_00000000100000000000000000000000};
        bins mhpmcounter24_enabled  = {44'b110000011000_00000001000000000000000000000000};
        bins mhpmcounter25_enabled  = {44'b110000011001_00000010000000000000000000000000};
        bins mhpmcounter26_enabled  = {44'b110000011010_00000100000000000000000000000000};
        bins mhpmcounter27_enabled  = {44'b110000011011_00001000000000000000000000000000};
        bins mhpmcounter28_enabled  = {44'b110000011100_00010000000000000000000000000000};
        bins mhpmcounter29_enabled  = {44'b110000011101_00100000000000000000000000000000};
        bins mhpmcounter30_enabled  = {44'b110000011110_01000000000000000000000000000000};
        bins mhpmcounter31_enabled  = {44'b110000011111_10000000000000000000000000000000};

        bins cycle_disabled         = {44'b110000000000_11111111111111111111111111111110};
        bins time_disabled          = {44'b110000000001_11111111111111111111111111111101};
        bins instret_disabled       = {44'b110000000010_11111111111111111111111111111011};
        bins mhpmcounter3_disabled   = {44'b110000000011_11111111111111111111111111110111};
        bins mhpmcounter4_disabled   = {44'b110000000100_11111111111111111111111111101111};
        bins mhpmcounter5_disabled   = {44'b110000000101_11111111111111111111111111011111};
        bins mhpmcounter6_disabled   = {44'b110000000110_11111111111111111111111110111111};
        bins mhpmcounter7_disabled   = {44'b110000000111_11111111111111111111111101111111};
        bins mhpmcounter8_disabled   = {44'b110000001000_11111111111111111111111011111111};
        bins mhpmcounter9_disabled   = {44'b110000001001_11111111111111111111110111111111};
        bins mhpmcounter10_disabled  = {44'b110000001010_11111111111111111111101111111111};
        bins mhpmcounter11_disabled  = {44'b110000001011_11111111111111111111011111111111};
        bins mhpmcounter12_disabled  = {44'b110000001100_11111111111111111110111111111111};
        bins mhpmcounter13_disabled  = {44'b110000001101_11111111111111111101111111111111};
        bins mhpmcounter14_disabled  = {44'b110000001110_11111111111111111011111111111111};
        bins mhpmcounter15_disabled  = {44'b110000001111_11111111111111110111111111111111};
        bins mhpmcounter16_disabled  = {44'b110000010000_11111111111111101111111111111111};
        bins mhpmcounter17_disabled  = {44'b110000010001_11111111111111011111111111111111};
        bins mhpmcounter18_disabled  = {44'b110000010010_11111111111110111111111111111111};
        bins mhpmcounter19_disabled  = {44'b110000010011_11111111111101111111111111111111};
        bins mhpmcounter20_disabled  = {44'b110000010100_11111111111011111111111111111111};
        bins mhpmcounter21_disabled  = {44'b110000010101_11111111110111111111111111111111};
        bins mmhpmcounter22_disabled  = {44'b110000010110_11111111101111111111111111111111};
        bins mhpmcounter23_disabled  = {44'b110000010111_11111111011111111111111111111111};
        bins mhpmcounter24_disabled  = {44'b110000011000_11111110111111111111111111111111};
        bins mhpmcounter25_disabled  = {44'b110000011001_11111101111111111111111111111111};
        bins mhpmcounter26_disabled  = {44'b110000011010_11111011111111111111111111111111};
        bins mhpmcounter27_disabled  = {44'b110000011011_11110111111111111111111111111111};
        bins mhpmcounter28_disabled  = {44'b110000011100_11101111111111111111111111111111};
        bins mhpmcounter29_disabled  = {44'b110000011101_11011111111111111111111111111111};
        bins mhpmcounter30_disabled  = {44'b110000011110_10111111111111111111111111111111};
        bins mhpmcounter31_disabled  = {44'b110000011111_01111111111111111111111111111111};
}
        `ifdef XLEN32
        cp_hpmh_counth: coverpoint {ins.current.insn[31:20], ins.current.csr[12'hB03][31:0] } {
            bins cycleh_enabled         = {44'b110010000000_00000000000000000000000000000001};
            bins timeh_enabled          = {44'b110010000001_00000000000000000000000000000010};
            bins instreth_enabled       = {44'b110010000010_00000000000000000000000000000100};
            bins mhpmcounter3h_enabled   = {44'b110010000011_00000000000000000000000000001000};
            bins mhpmcounter4h_enabled   = {44'b110010000100_00000000000000000000000000010000};
            bins mpmcounter5h_enabled   = {44'b110010000101_00000000000000000000000000100000};
            bins mpmcounter6h_enabled   = {44'b110010000110_00000000000000000000000001000000};
            bins mhpmcounter7h_enabled   = {44'b110010000111_00000000000000000000000010000000};
            bins mhpmcounter8h_enabled   = {44'b110010001000_00000000000000000000000100000000};
            bins mhpmcounter9h_enabled   = {44'b110010001001_00000000000000000000001000000000};
            bins mhpmcounter10h_enabled  = {44'b110010001010_00000000000000000000010000000000};
            bins mhpmcounter11h_enabled  = {44'b110010001011_00000000000000000000100000000000};
            bins mhpmcounter12h_enabled  = {44'b110010001100_00000000000000000001000000000000};
            bins mhpmcounter13h_enabled  = {44'b110010001101_00000000000000000010000000000000};
            bins mhpmcounter14h_enabled  = {44'b110010001110_00000000000000000100000000000000};
            bins mhpmcounter15h_enabled  = {44'b110010001111_00000000000000001000000000000000};
            bins mhpmcounter16h_enabled  = {44'b110010010000_00000000000000010000000000000000};
            bins mhpmcounter17h_enabled  = {44'b110010010001_00000000000000100000000000000000};
            bins mhpmcounter18h_enabled  = {44'b110010010010_00000000000001000000000000000000};
            bins mhpmcounter19h_enabled  = {44'b110010010011_00000000000010000000000000000000};
            bins mhpmcounter20h_enabled  = {44'b110010010100_00000000000100000000000000000000};
            bins mhpmcounter21h_enabled  = {44'b110010010101_00000000001000000000000000000000};
            bins mhpmcounter22h_enabled  = {44'b110010010110_00000000010000000000000000000000};
            bins mhpmcounter23h_enabled  = {44'b110010010111_00000000100000000000000000000000};
            bins mhpmcounter24h_enabled  = {44'b110010011000_00000001000000000000000000000000};
            bins mhpmcounter25h_enabled  = {44'b110010011001_00000010000000000000000000000000};
            bins mhpmcounter26h_enabled  = {44'b110010011010_00000100000000000000000000000000};
            bins mhpmcounter27h_enabled  = {44'b110010011011_00001000000000000000000000000000};
            bins mhpmcounter28h_enabled  = {44'b110010011100_00010000000000000000000000000000};
            bins mmhpmcounter29h_enabled  = {44'b110010011101_00100000000000000000000000000000};
            bins mhpmcounter30h_enabled  = {44'b110010011110_01000000000000000000000000000000};
            bins mhpmcounter31h_enabled  = {44'b110010011111_10000000000000000000000000000000};

            bins cycleh_disabled         = {44'b110010000000_11111111111111111111111111111110};
            bins timeh_disabled          = {44'b110010000001_11111111111111111111111111111101};
            bins instreth_disabled       = {44'b110010000010_11111111111111111111111111111011};
            bins mhpmcounter3h_disabled   = {44'b110010000011_11111111111111111111111111110111};
            bins mhpmcounter4h_disabled   = {44'b110010000100_11111111111111111111111111101111};
            bins mhpmcounter5h_disabled   = {44'b110010000101_11111111111111111111111111011111};
            bins mhpmcounter6h_disabled   = {44'b110010000110_11111111111111111111111110111111};
            bins mhpmcounter7h_disabled   = {44'b110010000111_11111111111111111111111101111111};
            bins mhpmcounter8h_disabled   = {44'b110010001000_11111111111111111111111011111111};
            bins mhpmcounter9h_disabled   = {44'b110010001001_11111111111111111111110111111111};
            bins mhpmcounter10h_disabled  = {44'b110010001010_11111111111111111111101111111111};
            bins mhpmcounter11h_disabled  = {44'b110010001011_11111111111111111111011111111111};
            bins mhpmcounter12h_disabled  = {44'b110010001100_11111111111111111110111111111111};
            bins mhpmcounter13h_disabled  = {44'b110010001101_11111111111111111101111111111111};
            bins mhpmcounter14h_disabled  = {44'b110010001110_11111111111111111011111111111111};
            bins mhpmcounter15h_disabled  = {44'b110010001111_11111111111111110111111111111111};
            bins mhpmcounter16h_disabled  = {44'b110010010000_11111111111111101111111111111111};
            bins mhpmcounter17h_disabled  = {44'b110010010001_11111111111111011111111111111111};
            bins mhpmcounter18h_disabled  = {44'b110010010010_11111111111110111111111111111111};
            bins mhpmcounter19h_disabled  = {44'b110010010011_11111111111101111111111111111111};
            bins mhpmcounter20h_disabled  = {44'b110010010100_11111111111011111111111111111111};
            bins mhpmcounter21h_disabled  = {44'b110010010101_11111111110111111111111111111111};
            bins mhpmcounter22h_disabled  = {44'b110010010110_11111111101111111111111111111111};
            bins mhpmcounter23h_disabled  = {44'b110010010111_11111111011111111111111111111111};
            bins mhpmcounter24h_disabled  = {44'b110010011000_11111110111111111111111111111111};
            bins mhpmcounter25h_disabled  = {44'b110010011001_11111101111111111111111111111111};
            bins mhpmcounter26h_disabled  = {44'b110010011010_11111011111111111111111111111111};
            bins mhpmcounter27h_disabled  = {44'b110010011011_11110111111111111111111111111111};
            bins mhpmcounter28h_disabled  = {44'b110010011100_11101111111111111111111111111111};
            bins mhpmcounter29h_disabled  = {44'b110010011101_11011111111111111111111111111111};
            bins mhpmcounter30h_disabled  = {44'b110010011110_10111111111111111111111111111111};
            bins mhpmcounter31h_disabled  = {44'b110010011111_01111111111111111111111111111111};
        `endif
    }

    cp_hmp_write: cross cp_hpmh_count, priv_mode_m;

    `ifdef XLEN32  
        cp_hpmh_write: cross cp_hpmh_counth, priv_mode_m;
    `endif

function void zihpm_sample(int hart, int issue, ins_t ins);
    Zihpm_cg.sample(ins);
endfunction