///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
///////////////////////////////////////////

   EndianH_endian_cg = new();         EndianH_endian_cg.set_inst_name("obj_EndianH_endian");