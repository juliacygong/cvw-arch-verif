///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
///////////////////////////////////////////

    SvinvalH_cg = new(); SvinvalH_cg.set_inst_name("obj_SvinvalH");

    