///////////////////////////////////////////
//
// RISC-V Architectural Functional Coverage Covergroups Initialization File
//
///////////////////////////////////////////

    ZicntrH_mcounters_cg = new();         ZicntrH_mcounters_cg.set_inst_name("obj_hcounters");